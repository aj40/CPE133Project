`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Cal Poly SLO
// Engineer: Allison Lee and Alex Johnson
// 
// Create Date: 11/18/2020 10:26:32 AM
//////////////////////////////////////////////////////////////////////////////////


module stopwatch(
    input clk,
    input start_stop,
    input reset,
    output Seg,
    output decimal
    );
endmodule
